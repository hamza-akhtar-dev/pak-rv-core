`ifndef RISCV_SVH

`define RISCV_SVH

    `define OPCODE_RTYPE 7'b0110011
    `define OPCODE_ITYPE 7'b0010011
    `define OPCODE_STYPE 7'b0100011
    `define OPCODE_BTYPE 7'b1100011
    `define OPCODE_UTYPE 7'b0010111
    `define OPCODE_JTYPE 7'b1101111
    
`endif
